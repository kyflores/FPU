module fpu(input[31:0] opA, input[31:0] opB, output[55:0] result,)